module message (
    input [9:0] sx, sy,
    input data_en,
    output logic [2:0] paint_rgb
    );

    localparam TEXT_COLOR = 3'b110;
    localparam BACKGROUND_COLOR = 3'b001;

    localparam bit [0:14][0:19] HELLO_WORLD_BMAP = {
        20'b1010_1110_1000_1000_0110,
        20'b1010_1000_1000_1000_1010,
        20'b1110_1100_1000_1000_1010,
        20'b1010_1000_1000_1000_1010,
        20'b1010_1110_1110_1110_1100,
        20'b0000_0000_0000_0000_0000,
        20'b1010_0110_1110_1000_1100,
        20'b1010_1010_1010_1000_1010,
        20'b1010_1010_1100_1000_1010,
        20'b1110_1010_1010_1000_1010,
        20'b1110_1100_1010_1110_1110,
        20'b0000_0000_0000_0000_0000,
        20'b0000_0000_0000_0000_0000,
        20'b0000_0000_0000_0000_0000,
        20'b0000_0000_0000_0000_0000
    };
    localparam bit [0:14][0:19] HER_BMAP = {
        20'b1010_1110_1110_0000_0000,
        20'b1010_1000_1010_0000_0000,
        20'b0100_1100_1110_0000_0000,
        20'b1010_1000_1000_0000_0000,
        20'b1010_1110_1000_0000_0000,
        20'b0000_0000_0000_0000_0000,
        20'b1110_1010_1110_1000_1000,
        20'b1010_1010_1010_1000_1000,
        20'b1010_1110_1010_1100_1000,
        20'b1010_0010_1010_1010_1000,
        20'b1010_1110_1010_1100_1000,
        20'b0000_0000_0000_0000_0000,
        20'b0000_0000_0000_0000_0000,
        20'b0000_0000_0000_0000_0000,
        20'b0000_0000_0000_0000_0000
    };
    // bitmap: MSB first, so we can write pixels left to right
    //logic [0:19] bmap [15];  // 20 pixels by 15 lines
    //initial begin
     //   bmap[0]  = 20'b1010_1110_1000_1000_0110;
     //   bmap[1]  = 20'b1010_1000_1000_1000_1010;
    //    bmap[2]  = 20'b1110_1100_1000_1000_1010;
     //   bmap[3]  = 20'b1010_1000_1000_1000_1010;
    //    bmap[4]  = 20'b1010_1110_1110_1110_1100;
     //   bmap[5]  = 20'b0000_0000_0000_0000_0000;
    //    bmap[6]  = 20'b1010_0110_1110_1000_1100;
   //     bmap[7]  = 20'b1010_1010_1010_1000_1010;
   //     bmap[8]  = 20'b1010_1010_1100_1000_1010;
   //     bmap[9]  = 20'b1110_1010_1010_1000_1010;
   //     bmap[10] = 20'b1110_1100_1010_1110_1110;
   //     bmap[11] = 20'b0000_0000_0000_0000_0000;
   //     bmap[12] = 20'b0000_0000_0000_0000_0000;
   //     bmap[13] = 20'b0000_0000_0000_0000_0000;
   //     bmap[14] = 20'b0000_0000_0000_0000_0000;
   // end

    // paint at 32x scale in active screen area
    logic msg_place;
    logic [4:0] x;  // 20 columns need five bits
    logic [3:0] y;  // 15 rows need four bits
    always_comb begin
        x = sx[9:5];    // every 32 horizontal pixels
        y = sy[8:5];    // every 32 vertical pixels
        msg_place = (data_en) ? HER_BMAP[y][x]: 0;
    end
    
    assign paint_rgb = (msg_place) ? TEXT_COLOR : BACKGROUND_COLOR;
endmodule
